`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   22:22:33 12/15/2020
// Design Name:   mips
// Module Name:   E:/Project/Verilog/piplineForClassTest/testMips.v
// Project Name:  piplineForClassTest
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: mips
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module testMips;

	// Inputs
	reg clk;
	reg reset;
	reg interrupt;
	wire [31:0] addr;
	// Instantiate the Unit Under Test (UUT)
	mips uut (
		.clk(clk), 
		.reset(reset),
		.interrupt(interrupt),
		.addr(addr)
	);

	initial begin
		// Initialize Inputs
		clk = 0;
		reset = 1;
		interrupt = 0;
		// Wait 100 ns for global reset to finish
		#10;
        
		// Add stimulus here
		reset = 0;
		#10;
		// interrupt = 1;

	end
    always #5 clk = ~clk;
endmodule

